localparam		ETH_ADDR 	= 0;
localparam		ETH_LEN 	= 1;
localparam		ETH_ST   	= 2;

localparam		UART_ADDR 	= 3;
localparam		UART_LEN 	= 4;
localparam		UART_ST   	= 5;


localparam		SRC_IP 		= 50;
localparam		SRC_MAC_H 	= 51;
localparam		SRC_MAC_L 	= 52;
localparam		DES_IP 		= 53;
localparam		DES_MAC_H 	= 54;
localparam		DES_MAC_L 	= 55;
