
module PISO 
#( // INPUT PARAMETERS
    parameter DATA_IN_WIDTH  = 64,
    parameter DATA_OUT_WIDTH = 16
)( // PORTS
    input  wire                         CLK,
    input  wire                         RESET_N,
    input  wire                         ENABLE,
    input  wire [DATA_IN_WIDTH -1 : 0]  DATA_IN,
    output wire                         READY,
    output wire [DATA_OUT_WIDTH -1 : 0] DATA_OUT,
    output wire                         OUT_VALID,
    input  wire                         OUT_READY     
);

// ******************************************************************
// LOCALPARAMS
// ******************************************************************
    localparam integer NUM_SHIFTS = DATA_IN_WIDTH / DATA_OUT_WIDTH;
// ******************************************************************

// ******************************************************************
// WIRES and REGS
// ******************************************************************
  reg [NUM_SHIFTS -1    : 0]  shift_count;
  reg [DATA_IN_WIDTH -1 : 0]  serial;
// ******************************************************************

  assign OUT_VALID = |shift_count;
  assign READY = !(OUT_VALID);

  assign DATA_OUT = serial [DATA_OUT_WIDTH-1:0];

  always @(posedge CLK or negedge RESET_N)
  begin: SHIFTER_COUNT
    if (!RESET_N)
      shift_count <= 0;
    else if (ENABLE & READY)
      shift_count <= {shift_count[NUM_SHIFTS-2:0], 1'b1};
    else if (OUT_VALID & OUT_READY) 
      shift_count <= {shift_count[NUM_SHIFTS-2:0], 1'b0};
  end


always @(posedge CLK or negedge RESET_N)
begin: DATA_SHIFT
    if (!RESET_N)
        serial <= 0;
    else begin
        if (ENABLE & READY)
            serial <= DATA_IN;
        else if (OUT_VALID & OUT_READY)
            serial <= {{DATA_OUT_WIDTH{1'b0}}, serial[DATA_IN_WIDTH-1:DATA_OUT_WIDTH]};
    end
end


endmodule
