// This is a simple example.
// You can make a your own header file and set its path to settings.
// (Preferences > Package Settings > Verilog Gadget > Settings - User)
//
//      "header": "Packages/Verilog Gadget/template/verilog_header.v"
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2020 All rights reserved
// -----------------------------------------------------------------------------
// Author : zhouchch@pku.edu.cn
// File   : CCU.v
// Create : 2020-07-14 21:09:52
// Revise : 2020-08-13 10:33:19
// -----------------------------------------------------------------------------
module EDC #(
    parameter CRD_WIDTH         = 16,
    parameter CRD_DIM           = 3 
    )(
    input       [CRD_DIM    -1 : 0][CRD_WIDTH           -1 : 0] Crd0,
    input       [CRD_DIM    -1 : 0][CRD_WIDTH           -1 : 0] Crd1,
    output reg signed[CRD_WIDTH*2+$clog2(CRD_DIM)            -1 : 0] DistSqr
);
//=====================================================================================================================
// Constant Definition :
//=====================================================================================================================


//=====================================================================================================================
// Variable Definition :
//=====================================================================================================================


//=====================================================================================================================
// Logic Design 1: FSM
//=====================================================================================================================
integer  i;
reg signed [CRD_WIDTH + 1           -1 : 0] Diff;

always @(*) begin
    DistSqr = 0;
    Diff    = 0;
    for(i = 0; i < CRD_DIM; i = i + 1) begin
        Diff = {Crd0[i][CRD_WIDTH -1], $signed(Crd0[i])} - {Crd1[i][CRD_WIDTH -1], $signed(Crd1[i])};
        DistSqr = DistSqr + Diff*Diff;
    end
end


//=====================================================================================================================
// Sub-Module :
//=====================================================================================================================



endmodule
