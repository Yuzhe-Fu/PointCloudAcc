module CTR #(
    parameters
) (
    ports
);
    
endmodule