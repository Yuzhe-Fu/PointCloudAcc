//-----------------------------------------------------------
//Simple Log2 calculation function
//-----------------------------------------------------------

`define CEIL(a,b) ( \
 (a%b)? (a/b+1):(a/b) \
)